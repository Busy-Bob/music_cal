module key_out(input IN_clk, input [3:0] IN_value, input IN_key, 
               output reg [3:0] OUT_col, output reg [7:0] OUT_SRCH, output reg [7:0] OUT_SRCL, output reg [7:0] OUT_DSTH, output reg [7:0] OUT_DSTL, output reg [3:0] OUT_ALU_OP, output reg OUT_finish);

endmodule 