library verilog;
use verilog.vl_types.all;
entity key_out_vlg_tst is
end key_out_vlg_tst;
