library verilog;
use verilog.vl_types.all;
entity debug_vlg_tst is
end debug_vlg_tst;
